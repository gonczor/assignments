library verilog;
use verilog.vl_types.all;
entity tester_vlg_vec_tst is
end tester_vlg_vec_tst;
