library verilog;
use verilog.vl_types.all;
entity Eight_Bit_Counter_vlg_vec_tst is
end Eight_Bit_Counter_vlg_vec_tst;
