library verilog;
use verilog.vl_types.all;
entity D_vhdl_vlg_sample_tst is
    port(
        KEY             : in     vl_logic_vector(0 downto 0);
        sampler_tx      : out    vl_logic
    );
end D_vhdl_vlg_sample_tst;
