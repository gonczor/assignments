library verilog;
use verilog.vl_types.all;
entity D_vhdl_vlg_vec_tst is
end D_vhdl_vlg_vec_tst;
